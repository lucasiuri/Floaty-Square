pll3M9Hz_inst : pll3M9Hz PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
