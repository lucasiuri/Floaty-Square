divFreq60Hz_inst : divFreq60Hz PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
